/*****************************************************************************
 *                                                                           *
 * Module:       Lab4                                                       *
 * Description:                                                              *
 *      This module is the top level module of MT3TB4 Lab 4                    *
 *                                                                           *
 *****************************************************************************/

module lab4 (
input				CLOCK_50,	
input		[0:0]	KEY, 
input 	[7:0] SW,               //for reset
output 	[7:0] LEDR,

// Bidirectionals
inout		[15:0]		DRAM_DQ,

// Outputs

output		[12:0]	DRAM_ADDR,
output 		[1:0]		DRAM_BA,
output					DRAM_LDQM,  //data mask; when it is low, the DQ is valid for reading and writing. 
output					DRAM_UDQM,
output					DRAM_RAS_N,
output 					DRAM_CAS_N,
output 					DRAM_CLK,
output					DRAM_CKE,
output 					DRAM_WE_N,
output 					DRAM_CS_N


);


// Internal Wires
wire [31:0] address;
wire bus_enable;
wire [1:0] byte_enable;
wire [15:0] write_data;
wire [15:0] read_data;
wire rw;
wire acknowledge;
wire SRAM_CE_N_wire;
wire SRAM_WE_N_wire;
wire SRAM_OE_N_wire;
wire SRAM_UB_N_wire;
wire SRAM_LB_N_wire;
assign SRAM_CE_N = SRAM_CE_N_wire;
assign SRAM_WE_N = SRAM_WE_N_wire;
assign SRAM_OE_N = SRAM_OE_N_wire;
assign SRAM_UB_N = SRAM_UB_N_wire;
assign SRAM_LB_N = SRAM_LB_N_wire;



assign LEDR=SW;

//Instantiate your sopc_system module generated by Platform Designer.  


sopc_system  controller (
		// example ports 
		.clk_clk(CLOCK_50),              
		.reset_reset_n(KEY[0]),        
		.sdram_clk_clk(DRAM_CLK),
		// more ports
		.sdram_addr_export(DRAM_ADDR),  
		.sdram_ba_export(DRAM_BA),    
		.sdram_cas_n_export(DRAM_CAS_N), 
		.sdram_cke_export(DRAM_CKE),   
		.sdram_cs_n_export(DRAM_CS_N),  
		.sdram_dq_export(DRAM_DQ),    
		.sdram_ldaqm_export(DRAM_LDQM),  
		.sdram_ras_n_export(DRAM_RAS_N), 
		.sdram_udqm_export(DRAM_UDQM),  
		.sdram_we_n_export(DRAM_WE_N),
		/*
		.sram_controller_0_conduit_end_export(SRAM_DQ), 
		.sram_controller_0_conduit_end_1_export(SRAM_ADDR), 
		.sram_controller_0_conduit_end_2_export(SRAM_CE_N_wire), 
		.sram_controller_0_conduit_end_3_export(SRAM_WE_N_wire), 
		.sram_controller_0_conduit_end_4_export(SRAM_OE_N_wire), 
		.sram_controller_0_conduit_end_5_export(SRAM_UB_N_wire), 
		.sram_controller_0_conduit_end_6_export(SRAM_LB_N_wire), 
		*/
	);

	
	

	
endmodule